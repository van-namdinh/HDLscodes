library verilog;
use verilog.vl_types.all;
entity seq_TLAT_X1 is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end seq_TLAT_X1;
