/*
 * Project name   :
 * File name      : 01Wire.v
 * Created date   : Th08 17 2018
 * Author         : Van-Nam DINH 
 * Last modified  : Th08 17 2018 09:05
 * Desc           :
 */
/*
#Link ref for doing this task
http://hdlbits.01xz.net/wiki/Exams/m2014_q4h
*/
module top_module(
    input   in,
    output  out);
    assign out = in;
endmodule
