/*
 * Project name   :
 * File name      : Wire4.v
 * Created date   : Th08 17 2018
 * Author         : Van-Nam DINH 
 * Last modified  : Th08 17 2018 14:23
 * Desc           :
 */

module top_module(
    input a,b,c,
    output  w,x,y,z);
assign w = a;
assign x = b;
assign y = b;
assign z = c;
endmodule

